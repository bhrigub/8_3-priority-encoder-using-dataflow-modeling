library verilog;
use verilog.vl_types.all;
entity tenco_p is
end tenco_p;
